magic
tech sky130A
magscale 1 2
timestamp 1729247295
<< nwell >>
rect -24 -1129 1868 140
<< nsubdiff >>
rect 12 70 72 104
rect 1772 70 1832 104
rect 12 44 46 70
rect 1798 44 1832 70
rect 12 -1059 46 -1033
rect 1798 -1059 1832 -1033
rect 12 -1093 72 -1059
rect 1772 -1093 1832 -1059
<< nsubdiffcont >>
rect 72 70 1772 104
rect 12 -1033 46 44
rect 1798 -1033 1832 44
rect 72 -1093 1772 -1059
<< poly >>
rect 201 -63 267 -47
rect 201 -97 217 -63
rect 251 -97 267 -63
rect 201 -113 267 -97
rect 1571 -64 1637 -48
rect 1571 -98 1587 -64
rect 1621 -98 1637 -64
rect 218 -136 248 -113
rect 1571 -114 1637 -98
rect 1589 -130 1619 -114
rect 218 -869 248 -854
rect 1589 -869 1619 -845
rect 200 -885 266 -869
rect 200 -919 216 -885
rect 250 -919 266 -885
rect 200 -935 266 -919
rect 1571 -885 1637 -869
rect 1571 -919 1587 -885
rect 1621 -919 1637 -885
rect 1571 -935 1637 -919
<< polycont >>
rect 217 -97 251 -63
rect 1587 -98 1621 -64
rect 216 -919 250 -885
rect 1587 -919 1621 -885
<< locali >>
rect 12 70 72 104
rect 1772 70 1832 104
rect 12 44 46 70
rect 1798 44 1832 70
rect 172 -97 217 -63
rect 251 -97 294 -63
rect 172 -149 206 -97
rect 260 -149 294 -97
rect 1543 -98 1587 -64
rect 1621 -98 1665 -64
rect 1543 -149 1577 -98
rect 1631 -149 1665 -98
rect 172 -885 206 -839
rect 260 -885 294 -839
rect 172 -919 216 -885
rect 250 -919 294 -885
rect 1543 -885 1577 -832
rect 1631 -885 1665 -832
rect 1543 -919 1587 -885
rect 1621 -919 1665 -885
rect 12 -1059 46 -1033
rect 1798 -1059 1832 -1033
rect 12 -1093 72 -1059
rect 1772 -1093 1832 -1059
<< viali >>
rect 217 -97 251 -63
rect 1587 -98 1621 -64
rect 216 -919 250 -885
rect 1587 -919 1621 -885
<< metal1 >>
rect 76 -22 525 40
rect 76 -956 138 -22
rect 205 -63 263 -57
rect 172 -97 217 -63
rect 251 -97 294 -63
rect 172 -103 294 -97
rect 172 -157 206 -103
rect 260 -150 294 -103
rect 449 -109 525 -22
rect 1313 -22 1761 40
rect 739 -112 749 -60
rect 801 -112 811 -60
rect 1027 -112 1037 -60
rect 1089 -112 1099 -60
rect 1313 -109 1389 -22
rect 1575 -64 1633 -58
rect 1543 -98 1587 -64
rect 1621 -98 1665 -64
rect 1543 -104 1665 -98
rect 1543 -150 1577 -104
rect 254 -162 385 -150
rect 254 -338 317 -162
rect 369 -338 385 -162
rect 254 -350 385 -338
rect 543 -350 719 -150
rect 831 -162 1007 -150
rect 831 -338 893 -162
rect 945 -338 1007 -162
rect 831 -350 1007 -338
rect 1119 -350 1295 -150
rect 1407 -162 1583 -150
rect 1631 -152 1665 -104
rect 1407 -332 1469 -162
rect 1452 -338 1469 -332
rect 1521 -338 1583 -162
rect 1452 -350 1583 -338
rect 608 -471 655 -350
rect 1183 -471 1230 -350
rect 1313 -437 1406 -391
rect 608 -518 1230 -471
rect 608 -638 655 -518
rect 1183 -638 1230 -518
rect 254 -650 430 -638
rect 254 -826 317 -650
rect 369 -826 430 -650
rect 172 -879 206 -832
rect 254 -838 430 -826
rect 543 -838 719 -638
rect 877 -649 961 -638
rect 877 -826 892 -649
rect 944 -826 961 -649
rect 877 -838 961 -826
rect 1119 -838 1295 -638
rect 1408 -650 1584 -638
rect 1408 -826 1469 -650
rect 1521 -826 1584 -650
rect 1408 -838 1584 -826
rect 260 -879 294 -838
rect 172 -885 294 -879
rect 172 -919 216 -885
rect 250 -919 294 -885
rect 204 -925 262 -919
rect 451 -928 461 -876
rect 513 -928 523 -876
rect 737 -925 1101 -879
rect 881 -956 957 -925
rect 1315 -928 1325 -876
rect 1377 -928 1387 -876
rect 1543 -879 1577 -838
rect 1631 -879 1665 -832
rect 1543 -885 1665 -879
rect 1543 -919 1587 -885
rect 1621 -919 1665 -885
rect 1575 -925 1633 -919
rect 1699 -956 1761 -22
rect 76 -1018 1761 -956
<< via1 >>
rect 749 -112 801 -60
rect 1037 -112 1089 -60
rect 317 -338 369 -162
rect 893 -338 945 -162
rect 1469 -338 1521 -162
rect 317 -826 369 -650
rect 892 -826 944 -649
rect 1469 -826 1521 -650
rect 461 -928 513 -876
rect 1325 -928 1377 -876
<< metal2 >>
rect 76 -22 1761 40
rect 76 -956 138 -22
rect 881 -50 957 -22
rect 738 -60 1101 -50
rect 738 -112 749 -60
rect 801 -112 1037 -60
rect 1089 -112 1101 -60
rect 738 -123 1101 -112
rect 317 -162 369 -150
rect 317 -471 369 -338
rect 891 -161 947 -151
rect 891 -348 947 -338
rect 1469 -162 1521 -149
rect 1469 -471 1521 -338
rect 317 -518 1521 -471
rect 315 -649 371 -639
rect 315 -836 371 -826
rect 892 -649 944 -518
rect 892 -838 944 -826
rect 1467 -650 1523 -640
rect 1467 -836 1523 -826
rect 449 -876 525 -866
rect 449 -928 461 -876
rect 513 -928 525 -876
rect 449 -956 525 -928
rect 76 -1018 525 -956
rect 1313 -876 1389 -866
rect 1313 -928 1325 -876
rect 1377 -928 1389 -876
rect 1313 -956 1389 -928
rect 1699 -956 1761 -22
rect 1313 -1018 1761 -956
<< via2 >>
rect 891 -162 947 -161
rect 891 -338 893 -162
rect 893 -338 945 -162
rect 945 -338 947 -162
rect 315 -650 371 -649
rect 315 -826 317 -650
rect 317 -826 369 -650
rect 369 -826 371 -650
rect 1467 -826 1469 -650
rect 1469 -826 1521 -650
rect 1521 -826 1523 -650
<< metal3 >>
rect 881 -161 957 -150
rect 881 -338 891 -161
rect 947 -338 957 -161
rect 881 -464 957 -338
rect 305 -524 1533 -464
rect 305 -649 381 -524
rect 305 -826 315 -649
rect 371 -826 381 -649
rect 305 -838 381 -826
rect 1457 -650 1533 -524
rect 1457 -826 1467 -650
rect 1523 -826 1533 -650
rect 1457 -838 1533 -826
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_0
timestamp 1729240876
transform 1 0 233 0 1 -738
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_1
timestamp 1729240876
transform 1 0 233 0 1 -250
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_2
timestamp 1729240876
transform 1 0 1604 0 1 -250
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_3
timestamp 1729240876
transform 1 0 1604 0 1 -738
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_VGK97L  sky130_fd_pr__pfet_01v8_VGK97L_0
timestamp 1729240876
transform 1 0 775 0 1 -250
box -144 -200 144 200
use sky130_fd_pr__pfet_01v8_VGK97L  sky130_fd_pr__pfet_01v8_VGK97L_1
timestamp 1729240876
transform 1 0 1351 0 1 -738
box -144 -200 144 200
use sky130_fd_pr__pfet_01v8_VGK97L  sky130_fd_pr__pfet_01v8_VGK97L_2
timestamp 1729240876
transform 1 0 1063 0 1 -250
box -144 -200 144 200
use sky130_fd_pr__pfet_01v8_VGK97L  sky130_fd_pr__pfet_01v8_VGK97L_3
timestamp 1729240876
transform 1 0 1351 0 1 -250
box -144 -200 144 200
use sky130_fd_pr__pfet_01v8_VGK97L  sky130_fd_pr__pfet_01v8_VGK97L_4
timestamp 1729240876
transform 1 0 487 0 1 -250
box -144 -200 144 200
use sky130_fd_pr__pfet_01v8_VGK97L  sky130_fd_pr__pfet_01v8_VGK97L_5
timestamp 1729240876
transform 1 0 487 0 1 -738
box -144 -200 144 200
use sky130_fd_pr__pfet_01v8_VGK97L  sky130_fd_pr__pfet_01v8_VGK97L_6
timestamp 1729240876
transform 1 0 775 0 1 -738
box -144 -200 144 200
use sky130_fd_pr__pfet_01v8_VGK97L  sky130_fd_pr__pfet_01v8_VGK97L_7
timestamp 1729240876
transform 1 0 1063 0 1 -738
box -144 -200 144 200
<< labels >>
flabel via2 338 -742 338 -742 0 FreeSans 480 0 0 0 D6
port 0 nsew
flabel via1 341 -248 341 -248 0 FreeSans 480 0 0 0 OUT
port 1 nsew
flabel metal2 910 12 910 12 0 FreeSans 480 0 0 0 VIN
port 2 nsew
flabel metal1 918 -976 918 -976 0 FreeSans 480 0 0 0 VIP
port 3 nsew
flabel nsubdiffcont 905 91 905 91 0 FreeSans 480 0 0 0 VDD
port 4 nsew
flabel metal1 630 -260 630 -260 0 FreeSans 480 0 0 0 D5
port 5 nsew
<< end >>
