magic
tech sky130A
magscale 1 2
timestamp 1729227955
<< nmos >>
rect -80 -100 80 100
<< ndiff >>
rect -138 88 -80 100
rect -138 -88 -126 88
rect -92 -88 -80 88
rect -138 -100 -80 -88
rect 80 88 138 100
rect 80 -88 92 88
rect 126 -88 138 88
rect 80 -100 138 -88
<< ndiffc >>
rect -126 -88 -92 88
rect 92 -88 126 88
<< poly >>
rect -80 172 80 188
rect -80 138 -64 172
rect 64 138 80 172
rect -80 100 80 138
rect -80 -138 80 -100
rect -80 -172 -64 -138
rect 64 -172 80 -138
rect -80 -188 80 -172
<< polycont >>
rect -64 138 64 172
rect -64 -172 64 -138
<< locali >>
rect -80 138 -64 172
rect 64 138 80 172
rect -126 88 -92 104
rect -126 -104 -92 -88
rect 92 88 126 104
rect 92 -104 126 -88
rect -80 -172 -64 -138
rect 64 -172 80 -138
<< viali >>
rect -45 138 45 172
rect -126 -88 -92 88
rect 92 -88 126 88
rect -45 -172 45 -138
<< metal1 >>
rect -57 172 57 178
rect -57 138 -45 172
rect 45 138 57 172
rect -57 132 57 138
rect -132 88 -86 100
rect -132 -88 -126 88
rect -92 -88 -86 88
rect -132 -100 -86 -88
rect 86 88 132 100
rect 86 -88 92 88
rect 126 -88 132 88
rect 86 -100 132 -88
rect -57 -138 57 -132
rect -57 -172 -45 -138
rect 45 -172 57 -138
rect -57 -178 57 -172
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 0.8 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 70 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
