magic
tech sky130A
magscale 1 2
timestamp 1729273826
<< nwell >>
rect -1962 -506 -962 2498
rect -334 1162 1936 2499
<< viali >>
rect -692 2359 -634 2405
rect 592 2371 626 2405
rect -693 2243 -634 2291
rect -693 2120 -634 2169
rect -693 1990 -633 2040
rect -692 1858 -632 1908
rect -693 1735 -634 1783
rect -810 716 -752 762
rect 239 716 297 762
<< metal1 >>
rect -1032 2439 637 2477
rect -1032 2283 -986 2439
rect -704 2405 -622 2439
rect 582 2411 637 2439
rect -704 2359 -692 2405
rect -634 2359 -622 2405
rect 580 2405 638 2411
rect 580 2371 592 2405
rect 626 2371 638 2405
rect 580 2365 638 2371
rect -704 2353 -622 2359
rect -705 2291 -197 2297
rect -705 2243 -693 2291
rect -634 2243 -197 2291
rect -705 2237 -197 2243
rect -705 2171 -622 2175
rect -705 2119 -693 2171
rect -634 2119 -622 2171
rect -705 2114 -622 2119
rect -705 2043 -621 2046
rect -705 1987 -694 2043
rect -633 1987 -621 2043
rect -705 1984 -621 1987
rect -704 1911 -620 1914
rect -704 1855 -692 1911
rect -632 1855 -620 1911
rect -704 1852 -620 1855
rect -705 1783 -497 1789
rect -705 1735 -693 1783
rect -634 1735 -497 1783
rect -144 1771 -134 1823
rect -82 1820 -72 1823
rect -82 1773 345 1820
rect -82 1771 -72 1773
rect -705 1729 -497 1735
rect -547 1374 -497 1729
rect -548 885 -497 1374
rect -548 843 1128 885
rect -1145 765 -740 768
rect -1145 713 -810 765
rect -752 713 -740 765
rect -1145 710 -740 713
rect 5 664 62 843
rect 1069 827 1128 843
rect 227 765 309 768
rect 227 713 239 765
rect 297 761 309 765
rect 297 715 668 761
rect 297 713 309 715
rect 227 710 309 713
rect -30 623 62 664
rect -30 560 27 623
rect -1363 -430 -1304 -283
rect 615 -430 674 -280
rect -1363 -479 674 -430
<< via1 >>
rect -693 2169 -634 2171
rect -693 2120 -634 2169
rect -693 2119 -634 2120
rect -694 2040 -633 2043
rect -694 1990 -693 2040
rect -693 1990 -633 2040
rect -694 1987 -633 1990
rect -692 1908 -632 1911
rect -692 1858 -632 1908
rect -692 1855 -632 1858
rect -134 1771 -82 1823
rect -810 762 -752 765
rect -810 716 -752 762
rect -810 713 -752 716
rect 239 762 297 765
rect 239 716 297 762
rect 239 713 297 716
<< metal2 >>
rect -705 2171 -187 2181
rect -705 2119 -693 2171
rect -634 2119 -187 2171
rect -705 2109 -187 2119
rect -936 2043 -343 2053
rect -936 1987 -694 2043
rect -633 1987 -343 2043
rect -936 1977 -343 1987
rect -936 668 -885 1977
rect -704 1911 -423 1921
rect -704 1855 -692 1911
rect -632 1855 -423 1911
rect -704 1845 -423 1855
rect -475 1017 -423 1845
rect -394 1151 -343 1977
rect -136 1825 -80 1835
rect -136 1759 -80 1769
rect 580 1451 634 1505
rect 580 1151 635 1451
rect -394 1098 635 1151
rect -474 989 -423 1017
rect -474 938 1286 989
rect 1061 937 1286 938
rect -810 765 297 775
rect -752 713 239 765
rect -810 703 297 713
rect -936 615 -629 668
rect -680 347 -629 615
rect 1214 612 1286 937
<< via2 >>
rect -136 1823 -80 1825
rect -136 1771 -134 1823
rect -134 1771 -82 1823
rect -82 1771 -80 1823
rect -136 1769 -80 1771
<< metal3 >>
rect -234 1825 -70 1830
rect -234 1769 -136 1825
rect -80 1769 -70 1825
rect -234 1764 -70 1769
rect -234 1728 -172 1764
rect -1153 1664 -172 1728
rect -4 667 72 1516
rect -257 607 72 667
rect -257 306 -181 607
use nmoscs  nmoscs_0
timestamp 1729225079
transform 1 0 812 0 1 187
box -328 -589 1054 655
use nmosgn  nmosgn_0
timestamp 1729233841
transform 1 0 -742 0 1 348
box -118 -750 1164 244
use pmoscs  pmoscs_0
timestamp 1729158591
transform 1 0 -1785 0 1 -342
box -177 -90 823 2773
use pmosgn  pmosgn_0
timestamp 1729247295
transform 1 0 -310 0 1 2291
box -24 -1129 1868 140
<< labels >>
flabel viali -661 2380 -661 2380 0 FreeSans 480 0 0 0 VDD
port 0 nsew
flabel viali -660 2269 -660 2269 0 FreeSans 480 0 0 0 VIP
port 1 nsew
flabel via1 -665 2147 -665 2147 0 FreeSans 480 0 0 0 VIN
port 2 nsew
flabel via1 -665 2012 -665 2012 0 FreeSans 480 0 0 0 OUT
port 3 nsew
flabel via1 -663 1883 -663 1883 0 FreeSans 480 0 0 0 RS
port 4 nsew
flabel viali -664 1756 -664 1756 0 FreeSans 480 0 0 0 GND
port 5 nsew
<< end >>
