magic
tech sky130A
magscale 1 2
timestamp 1729233841
<< psubdiff >>
rect -118 204 -58 238
rect 1104 204 1164 238
rect -118 178 -84 204
rect 1130 178 1164 204
rect -118 -710 -84 -684
rect 1130 -710 1164 -684
rect -118 -744 -58 -710
rect 1104 -744 1164 -710
<< psubdiffcont >>
rect -58 204 1104 238
rect -118 -684 -84 178
rect 1130 -684 1164 178
rect -58 -744 1104 -710
<< poly >>
rect -34 154 58 170
rect -34 120 -18 154
rect 16 120 58 154
rect -34 104 58 120
rect 28 93 58 104
rect 988 154 1080 170
rect 988 120 1030 154
rect 1064 120 1080 154
rect 988 104 1080 120
rect 988 92 1018 104
rect 117 -302 930 -204
rect 28 -610 58 -598
rect -34 -626 58 -610
rect -34 -660 -18 -626
rect 16 -660 58 -626
rect -34 -676 58 -660
rect 988 -610 1018 -598
rect 988 -626 1080 -610
rect 988 -660 1030 -626
rect 1064 -660 1080 -626
rect 988 -676 1080 -660
<< polycont >>
rect -18 120 16 154
rect 1030 120 1064 154
rect -18 -660 16 -626
rect 1030 -660 1064 -626
<< locali >>
rect -118 204 -58 238
rect 1104 204 1164 238
rect -118 178 -84 204
rect 1130 178 1164 204
rect -18 154 16 170
rect -18 74 16 120
rect 1030 154 1064 170
rect 1030 82 1064 120
rect -18 -626 16 -589
rect -18 -676 16 -660
rect 1030 -626 1064 -587
rect 1030 -676 1064 -660
rect -118 -710 -84 -684
rect 1130 -710 1164 -684
rect -118 -744 -58 -710
rect 1104 -744 1164 -710
<< viali >>
rect 724 204 758 238
rect -18 120 16 154
rect 1030 120 1064 154
rect -18 -660 16 -626
rect 1030 -660 1064 -626
rect 288 -744 322 -710
<< metal1 >>
rect 712 238 770 244
rect 712 204 724 238
rect 758 204 770 238
rect 712 198 770 204
rect -24 154 22 166
rect -24 120 -18 154
rect 16 120 22 154
rect -24 82 22 120
rect -24 70 114 82
rect -24 -106 61 70
rect 113 -106 123 70
rect -24 -118 114 -106
rect 282 -231 328 82
rect 487 -106 497 70
rect 549 -106 559 70
rect 718 -231 764 198
rect 1024 154 1070 166
rect 1024 120 1030 154
rect 1064 120 1070 154
rect 1024 82 1070 120
rect 931 70 1070 82
rect 923 -106 933 70
rect 985 -106 1070 70
rect 931 -118 1070 -106
rect 282 -275 764 -231
rect 64 -356 253 -310
rect 64 -388 110 -356
rect -30 -400 116 -388
rect -30 -576 61 -400
rect 113 -576 123 -400
rect -30 -588 116 -576
rect -24 -626 22 -588
rect -24 -660 -18 -626
rect 16 -660 22 -626
rect -24 -672 22 -660
rect 282 -704 328 -275
rect 487 -576 497 -400
rect 549 -576 559 -400
rect 718 -588 764 -275
rect 793 -356 982 -311
rect 937 -388 982 -356
rect 930 -400 1076 -388
rect 923 -576 933 -400
rect 985 -576 1076 -400
rect 930 -588 1076 -576
rect 1024 -626 1070 -588
rect 1024 -660 1030 -626
rect 1064 -660 1070 -626
rect 1024 -672 1070 -660
rect 276 -710 334 -704
rect 276 -744 288 -710
rect 322 -744 334 -710
rect 276 -750 334 -744
<< via1 >>
rect 61 -106 113 70
rect 497 -106 549 70
rect 933 -106 985 70
rect 61 -576 113 -400
rect 497 -576 549 -400
rect 933 -576 985 -400
<< metal2 >>
rect 51 70 123 82
rect 51 -106 61 70
rect 113 -106 123 70
rect 51 -231 123 -106
rect 495 70 551 80
rect 495 -116 551 -106
rect 924 70 996 82
rect 924 -106 933 70
rect 985 -106 996 70
rect 924 -231 996 -106
rect 51 -275 996 -231
rect 59 -400 115 -390
rect 59 -586 115 -576
rect 487 -400 559 -275
rect 487 -576 497 -400
rect 549 -576 559 -400
rect 487 -588 559 -576
rect 931 -400 987 -390
rect 931 -586 987 -576
<< via2 >>
rect 495 -106 497 70
rect 497 -106 549 70
rect 549 -106 551 70
rect 59 -576 61 -400
rect 61 -576 113 -400
rect 113 -576 115 -400
rect 931 -576 933 -400
rect 933 -576 985 -400
rect 985 -576 987 -400
<< metal3 >>
rect 485 70 561 82
rect 485 -106 495 70
rect 551 -106 561 70
rect 485 -224 561 -106
rect 49 -284 997 -224
rect 49 -400 125 -284
rect 49 -576 59 -400
rect 115 -576 125 -400
rect 49 -588 125 -576
rect 921 -400 997 -284
rect 921 -576 931 -400
rect 987 -576 997 -400
rect 921 -588 997 -576
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_0
timestamp 1729227955
transform 1 0 43 0 1 -18
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_1
timestamp 1729227955
transform 1 0 1003 0 1 -18
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_2
timestamp 1729227955
transform 1 0 1003 0 1 -488
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_3
timestamp 1729227955
transform 1 0 43 0 1 -488
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_DXNGNZ  sky130_fd_pr__nfet_01v8_DXNGNZ_0
timestamp 1729227955
transform 1 0 523 0 1 -488
box -465 -188 465 188
use sky130_fd_pr__nfet_01v8_DXNGNZ  sky130_fd_pr__nfet_01v8_DXNGNZ_1
timestamp 1729227955
transform 1 0 523 0 1 -18
box -465 -188 465 188
<< labels >>
flabel via1 84 -16 84 -16 0 FreeSans 480 0 0 0 OUT
port 0 nsew
flabel via1 87 -493 87 -493 0 FreeSans 480 0 0 0 D6
port 1 nsew
flabel metal1 306 -494 306 -494 0 FreeSans 480 0 0 0 GND
port 2 nsew
<< end >>
