magic
tech sky130A
magscale 1 2
timestamp 1729158591
<< nwell >>
rect -177 -90 823 2773
<< nsubdiff >>
rect -141 2703 -81 2737
rect 727 2703 787 2737
rect -141 2677 -107 2703
rect 753 2677 787 2703
rect -141 -19 -107 7
rect 753 -19 787 7
rect -141 -53 -81 -19
rect 727 -53 787 -19
<< nsubdiffcont >>
rect -81 2703 727 2737
rect -141 7 -107 2677
rect 753 7 787 2677
rect -81 -53 727 -19
<< poly >>
rect -58 2665 36 2681
rect -58 2631 -42 2665
rect -8 2631 36 2665
rect -58 2615 36 2631
rect 6 2608 36 2615
rect 610 2665 704 2681
rect 610 2631 654 2665
rect 688 2631 704 2665
rect 610 2615 704 2631
rect 610 2608 640 2615
rect -58 1970 36 1986
rect 94 1984 294 2086
rect -58 1936 -42 1970
rect -8 1936 36 1970
rect -58 1920 36 1936
rect 6 1913 36 1920
rect 610 1971 704 1987
rect 610 1937 654 1971
rect 688 1937 704 1971
rect 610 1921 704 1937
rect 610 1914 640 1921
rect -58 1276 36 1292
rect 94 1290 552 1392
rect -58 1242 -42 1276
rect -8 1242 36 1276
rect -58 1226 36 1242
rect 6 1219 36 1226
rect 610 1277 704 1293
rect 610 1243 654 1277
rect 688 1243 704 1277
rect 610 1227 704 1243
rect 610 1220 640 1227
rect -58 583 36 599
rect 352 596 552 698
rect -58 549 -42 583
rect -8 549 36 583
rect -58 533 36 549
rect 6 526 36 533
rect 610 583 704 599
rect 610 549 654 583
rect 688 549 704 583
rect 610 533 704 549
rect 610 526 640 533
<< polycont >>
rect -42 2631 -8 2665
rect 654 2631 688 2665
rect -42 1936 -8 1970
rect 654 1937 688 1971
rect -42 1242 -8 1276
rect 654 1243 688 1277
rect -42 549 -8 583
rect 654 549 688 583
<< locali >>
rect -141 2703 -81 2737
rect 727 2703 787 2737
rect -141 2677 -107 2703
rect 753 2677 787 2703
rect -58 2631 -42 2665
rect -8 2631 8 2665
rect 638 2631 654 2665
rect 688 2631 704 2665
rect -40 2576 -6 2631
rect 652 2584 686 2631
rect -58 1936 -42 1970
rect -8 1936 8 1970
rect 638 1937 654 1971
rect 688 1937 704 1971
rect -40 1881 -6 1936
rect 652 1884 686 1937
rect -58 1242 -42 1276
rect -8 1242 8 1276
rect 638 1243 654 1277
rect 688 1243 704 1277
rect -40 1186 -6 1242
rect 652 1188 686 1243
rect -58 549 -42 583
rect -8 549 8 583
rect 638 549 654 583
rect 688 549 704 583
rect -40 501 -6 549
rect 652 502 686 549
rect -141 -19 -107 7
rect 753 -19 787 7
rect -141 -53 -81 -19
rect 727 -53 787 -19
<< viali >>
rect -42 2631 -8 2665
rect 654 2631 688 2665
rect 753 2631 787 2665
rect -42 1936 -8 1970
rect 654 1937 688 1971
rect -42 1242 -8 1276
rect 654 1243 688 1277
rect -141 549 -107 583
rect -42 549 -8 583
rect 654 549 688 583
<< metal1 >>
rect -54 2665 4 2671
rect -54 2631 -42 2665
rect -8 2631 4 2665
rect -54 2625 4 2631
rect 642 2665 799 2671
rect 642 2631 654 2665
rect 688 2631 753 2665
rect 787 2631 799 2665
rect 642 2625 799 2631
rect -46 2582 0 2625
rect 646 2582 692 2625
rect -52 2572 86 2582
rect -60 2194 -50 2572
rect 2 2194 86 2572
rect -52 2182 86 2194
rect 300 2144 346 2582
rect 558 2224 692 2582
rect 556 2182 692 2224
rect 556 2144 606 2182
rect 300 2092 606 2144
rect -54 1970 4 1976
rect -54 1936 -42 1970
rect -8 1936 4 1970
rect -54 1930 4 1936
rect -46 1884 0 1930
rect -45 1881 0 1884
rect -58 1500 -48 1876
rect 4 1500 38 1876
rect 92 1500 102 1876
rect -6 1490 44 1500
rect -54 1276 4 1282
rect -54 1242 -42 1276
rect -8 1242 4 1276
rect -54 1236 4 1242
rect -46 1194 0 1236
rect 40 1234 266 1280
rect 40 1194 90 1234
rect -46 794 90 1194
rect 300 590 346 2092
rect 642 1971 700 1977
rect 642 1937 654 1971
rect 688 1937 700 1971
rect 642 1931 700 1937
rect 646 1888 692 1931
rect 558 1488 692 1888
rect 558 1448 604 1488
rect 392 1402 604 1448
rect 642 1277 700 1283
rect 642 1243 654 1277
rect 688 1243 700 1277
rect 642 1237 700 1243
rect 646 1187 692 1237
rect 544 806 554 1182
rect 608 806 644 1182
rect 696 806 706 1182
rect -153 583 4 589
rect -153 549 -141 583
rect -107 549 -42 583
rect -8 549 4 583
rect -153 543 4 549
rect -46 500 0 543
rect 42 538 346 590
rect 642 583 700 589
rect 642 549 654 583
rect 688 549 700 583
rect 642 543 700 549
rect 42 500 88 538
rect -46 100 88 500
rect 300 100 346 538
rect 646 498 692 543
rect 602 490 646 492
rect 544 112 554 490
rect 606 488 646 490
rect 606 112 643 488
rect 695 112 705 488
rect 602 108 646 112
<< via1 >>
rect -50 2194 2 2572
rect -48 1500 4 1876
rect 38 1500 92 1876
rect 554 806 608 1182
rect 644 806 696 1182
rect 554 112 606 490
rect 643 112 695 488
<< metal2 >>
rect -52 2582 6 2592
rect -62 2182 -52 2582
rect 6 2182 86 2582
rect -52 2172 6 2182
rect 38 1888 104 1890
rect -52 1876 104 1888
rect -52 1500 -48 1876
rect 4 1500 38 1876
rect 92 1500 104 1876
rect -52 1488 104 1500
rect 26 1372 102 1488
rect 26 1314 620 1372
rect 544 1196 620 1314
rect 544 1182 698 1196
rect 544 806 554 1182
rect 608 806 644 1182
rect 696 806 698 1182
rect 544 794 698 806
rect 640 500 698 510
rect 552 492 608 500
rect 552 490 640 492
rect 608 112 640 490
rect 552 108 640 112
rect 552 102 608 108
rect 640 90 698 100
<< via2 >>
rect -52 2572 6 2582
rect -52 2194 -50 2572
rect -50 2194 2 2572
rect 2 2194 6 2572
rect -52 2182 6 2194
rect 552 112 554 490
rect 554 112 606 490
rect 606 112 608 490
rect 640 488 698 500
rect 640 112 643 488
rect 643 112 695 488
rect 695 112 698 488
rect 640 100 698 112
<< metal3 >>
rect -62 2582 86 2594
rect -62 2182 -52 2582
rect 6 2182 86 2582
rect -62 2170 86 2182
rect -62 2070 16 2170
rect -62 2006 708 2070
rect -62 674 16 2006
rect 630 1659 708 2006
rect 630 674 709 1659
rect -62 610 709 674
rect -62 609 16 610
rect 630 508 709 610
rect 540 500 709 508
rect 540 490 640 500
rect 540 112 552 490
rect 608 112 640 490
rect 540 100 640 112
rect 698 100 709 500
rect 540 90 709 100
rect 631 89 709 90
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_0
timestamp 1729132909
transform 1 0 625 0 1 1688
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_1
timestamp 1729132909
transform 1 0 21 0 1 300
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_2
timestamp 1729132909
transform 1 0 625 0 1 300
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_3
timestamp 1729132909
transform 1 0 21 0 1 994
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_4
timestamp 1729132909
transform 1 0 625 0 1 994
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_5
timestamp 1729132909
transform 1 0 21 0 1 1688
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_6
timestamp 1729132909
transform 1 0 625 0 1 2382
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_7
timestamp 1729132909
transform 1 0 21 0 1 2382
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_0
timestamp 1729150525
transform 1 0 323 0 1 2382
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_1
timestamp 1729150525
transform 1 0 323 0 1 1688
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_2
timestamp 1729150525
transform 1 0 323 0 1 994
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_3
timestamp 1729150525
transform 1 0 323 0 1 300
box -323 -300 323 300
<< labels >>
flabel metal1 722 2641 722 2641 0 FreeSans 160 0 0 0 VDD
port 0 nsew
flabel metal3 524 2035 530 2035 0 FreeSans 160 0 0 0 D5
port 1 nsew
flabel metal2 570 1327 570 1327 0 FreeSans 160 0 0 0 D1
port 2 nsew
flabel metal1 566 1436 566 1436 0 FreeSans 160 0 0 0 D2
port 3 nsew
<< end >>
